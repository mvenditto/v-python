module py_test
import py

#flag -L/usr/lib/python3.9/config-3.9-x86_64-linux-gnu 
#flag -L/usr/lib/x86_64-linux-gnu
#flag -lcrypt 
#flag -lpython3.9
#flag -ldl 
#flag -lm

fn testsuite_begin() {
	
}

fn testsuite_end() {
	
}
